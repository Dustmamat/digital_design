LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY TBLAB2ES1 IS
END TBLAB2ES1;
ARCHITECTURE BHV OF TBLAB2ES1 IS
	COMPONENT lab2part1
        PORT (
            SW: IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
            HEX0: OUT STD_LOGIC_VECTOR (6 DOWNTO 0));
	END COMPONENT;
SIGNAL C: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL DECOUT : STD_LOGIC_VECTOR (6 DOWNTO 0);
BEGIN
	DISPLAYOUT: lab2part1 PORT MAP (
        SW=>C,
        HEX0 => DECOUT);
	PROCESS
	BEGIN
	C(0)<='0';
	C(1)<='0';
	C(2)<='0';
	WAIT FOR 20 ns;

	C(2)<='1';
	WAIT FOR 20 ns;
	C(1)<='1';
	WAIT FOR 20 ns;
	C(2)<='0';
	WAIT FOR 20 ns;
	C(0)<='1';
	WAIT for 20 ns;
	WAIT;
	END PROCESS;

END BHV;