LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY mux2to1 IS 
	PORT(
	X: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	Y: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	S: IN STD_LOGIC;
	M: OUT STD_LOGIC_VECTOR (2 DOWNTO 0));
END ENTITY;

ARCHITECTURE STR OF MUX2TO1 IS
	BEGIN
	PROCESS (X, Y, S)
	BEGIN
	M(0)<=(NOT S AND X(0)) OR (S AND Y(0));
	M(1)<=(NOT S AND X(1)) OR (S AND Y(1));
	M(2)<=(NOT S AND X(2)) OR (S AND Y(2));
	END PROCESS;
END ARCHITECTURE;
	
